----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    22:58:06 09/17/2014 
-- Design Name: 
-- Module Name:    dev_select - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity dev_select is
PORT (a: in std_logic_vector(7 downto 0);
		y: out std_logic_vector(2 downto 0)
		);
end dev_select;

architecture Behavioral of dev_select is
begin

		---with a(7) select
		---y <= "111" when '1',
		----"000" when others;
		
		
		
		
	--y(2) <= (a(4) and not a(5) and not a(6) and not a(7)) or
---			(a(5) and not a(6) and not a(7)) or
			---(a(6) and not a(7)) or a(7);
			
	---y(1) <= (a(2) and not a(3) and not a(4) and not a(5) and not a(6) and not a(7)) or
			---(a(3) and not a(4) and not a(5) and not a(6) and not a(7)) or
			---(a(6) and not a(7)) or a(7);
			
	---y(0) <= (a(1) and not a(2) and not a(3) and not a(4) and not a(5) and not a(6) and not a(7)) or
			---(a(3) and not a(4) and not a(5) and not a(6) and not a(7)) or
			---(a(5) and not a(6) and not a(7)) or a(7);
			
	with a select
		y <= "000" when "00000001",
		"001" when "00000010",
		"001" when "00000011",
		"010" when "00000100",
		"010" when "00000101",
		"010" when "00000110",
		"010" when "00000111",
		"011" when "00001000",
		"011" when "00001001",
		"011" when "00001010",
		"011" when "00001011",
		"011" when "00001100",
		"011" when "00001101",
		"011" when "00001110",
		"011" when "00001111",
		"100" when "00010000",
		"100" when "00010001",
		"100" when "00010010",
		"100" when "00010011",
		"100" when "00010100",
		"100" when "00010101",
		"100" when "00010110",
		"100" when "00010111",
		"100" when "00011000",
		"100" when "00011001",
		"100" when "00011010",
		"100" when "00011011",
		"100" when "00011100",
		"100" when "00011101",
		"100" when "00011110",
		"100" when "00011111",
		"101" when "00100000",
		"101" when "00100001",
		"101" when "00100010",
		"101" when "00100011",
		"101" when "00100100",
		"101" when "00100101",
		"101" when "00100110",
		"101" when "00100111",
		"101" when "00101000",
		"101" when "00101001",
		"101" when "00101010",
		"101" when "00101011",
		"101" when "00101100",
		"101" when "00101101",
		"101" when "00101110",
		"101" when "00101111",
		"101" when "00110000",
		"101" when "00110001",
		"101" when "00110010",
		"101" when "00110011",
		"101" when "00110100",
		"101" when "00110101",
		"101" when "00110110",
		"101" when "00110111",
		"101" when "00111000",
		"101" when "00111001",
		"101" when "00111010",
		"101" when "00111011",
		"101" when "00111100",
		"101" when "00111101",
		"101" when "00111110",
		"101" when "00111111",
		"110" when "01000000",
		"110" when "01000001",
		"110" when "01000010",
		"110" when "01000011",
		"110" when "01000100",
		"110" when "01000101",
		"110" when "01000110",
		"110" when "01000111",
		"110" when "01001000",
		"110" when "01001001",
		"110" when "01001010",
		"110" when "01001011",
		"110" when "01001100",
		"110" when "01001101",
		"110" when "01001110",
		"110" when "01001111",
		"110" when "01010000",
		"110" when "01010001",
		"110" when "01010010",
		"110" when "01010011",
		"110" when "01010100",
		"110" when "01010101",
		"110" when "01010110",
		"110" when "01010111",
		"110" when "01011000",
		"110" when "01011001",
		"110" when "01011010",
		"110" when "01011011",
		"110" when "01011100",
		"110" when "01011101",
		"110" when "01011110",
		"110" when "01011111",
		"110" when "01100000",
		"110" when "01100001",
		"110" when "01100010",
		"110" when "01100011",
		"110" when "01100100",
		"110" when "01100101",
		"110" when "01100110",
		"110" when "01100111",
		"110" when "01101000",
		"110" when "01101001",
		"110" when "01101010",
		"110" when "01101011",
		"110" when "01101100",
		"110" when "01101101",
		"110" when "01101110",
		"110" when "01101111",
		"110" when "01110000",
		"110" when "01110001",
		"110" when "01110010",
		"110" when "01110011",
		"110" when "01110100",
		"110" when "01110101",
		"110" when "01110110",
		"110" when "01110111",
		"110" when "01111000",
		"110" when "01111001",
		"110" when "01111010",
		"110" when "01111011",
		"110" when "01111100",
		"110" when "01111101",
		"110" when "01111110",
		"110" when "01111111",
		"111" when "10000000",
		"111" when "10000001",
		"111" when "10000010",
		"111" when "10000011",
		"111" when "10000100",
		"111" when "10000101",
		"111" when "10000110",
		"111" when "10000111",
		"111" when "10001000",
		"111" when "10001001",
		"111" when "10001010",
		"111" when "10001011",
		"111" when "10001100",
		"111" when "10001101",
		"111" when "10001110",
		"111" when "10001111",
		"111" when "10010000",
		"111" when "10010001",
		"111" when "10010010",
		"111" when "10010011",
		"111" when "10010100",
		"111" when "10010101",
		"111" when "10010110",
		"111" when "10010111",
		"111" when "10011000",
		"111" when "10011001",
		"111" when "10011010",
		"111" when "10011011",
		"111" when "10011100",
		"111" when "10011101",
		"111" when "10011110",
		"111" when "10011111",
		"111" when "10100000",
		"111" when "10100001",
		"111" when "10100010",
		"111" when "10100011",
		"111" when "10100100",
		"111" when "10100101",
		"111" when "10100110",
		"111" when "10100111",
		"111" when "10101000",
		"111" when "10101001",
		"111" when "10101010",
		"111" when "10101011",
		"111" when "10101100",
		"111" when "10101101",
		"111" when "10101110",
		"111" when "10101111",
		"111" when "10110000",
		"111" when "10110001",
		"111" when "10110010",
		"111" when "10110011",
		"111" when "10110100",
		"111" when "10110101",
		"111" when "10110110",
		"111" when "10110111",
		"111" when "10111000",
		"111" when "10111001",
		"111" when "10111010",
		"111" when "10111011",
		"111" when "10111100",
		"111" when "10111101",
		"111" when "10111110",
		"111" when "10111111",
		"111" when "11000000",
		"111" when "11000001",
		"111" when "11000010",
		"111" when "11000011",
		"111" when "11000100",
		"111" when "11000101",
		"111" when "11000110",
		"111" when "11000111",
		"111" when "11001000",
		"111" when "11001001",
		"111" when "11001010",
		"111" when "11001011",
		"111" when "11001100",
		"111" when "11001101",
		"111" when "11001110",
		"111" when "11001111",
		"111" when "11010000",
		"111" when "11010001",
		"111" when "11010010",
		"111" when "11010011",
		"111" when "11010100",
		"111" when "11010101",
		"111" when "11010110",
		"111" when "11010111",
		"111" when "11011000",
		"111" when "11011001",
		"111" when "11011010",
		"111" when "11011011",
		"111" when "11011100",
		"111" when "11011101",
		"111" when "11011110",
		"111" when "11011111",
		"111" when "11100000",
		"111" when "11100001",
		"111" when "11100010",
		"111" when "11100011",
		"111" when "11100100",
		"111" when "11100101",
		"111" when "11100110",
		"111" when "11100111",
		"111" when "11101000",
		"111" when "11101001",
		"111" when "11101010",
		"111" when "11101011",
		"111" when "11101100",
		"111" when "11101101",
		"111" when "11101110",
		"111" when "11101111",
		"111" when "11110000",
		"111" when "11110001",
		"111" when "11110010",
		"111" when "11110011",
		"111" when "11110100",
		"111" when "11110101",
		"111" when "11110110",
		"111" when "11110111",
		"111" when "11111000",
		"111" when "11111001",
		"111" when "11111010",
		"111" when "11111011",
		"111" when "11111100",
		"111" when "11111101",
		"111" when "11111110",
		"111" when "11111111",
		"000" when others;
			
			

	
end Behavioral;

