package Common is    -- untested...

   type finit_state is (start, bit_0, bit_1, bit_2, bit_3, bit_4, bit_5, stop);

   -- (optional) useful tools

end Common;

package body Common is
   -- subprogram bodies here
end Common;